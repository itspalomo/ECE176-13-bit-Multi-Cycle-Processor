// this is a test

module test ():
    
endmodule
	
//////////////////////////////////////////////////////////////////////////////////
// Class: ECE 176
// Team Members: Jose Maciel Torres, Subham Savita
// 
// Design Name: Top Level Design Test Bench
// Module Name: risc_proc_tb
// Project Name: 13-bit RISC Processor
// Description: 
// 			
//				
// Port List: 
//			
//	
//////////////////////////////////////////////////////////////////////////////////
module risc_proc_tb();
	
endmodule
// this is a test

module test ():
wire [3:0] test1;    
endmodule